package weight_pkg;

  parameter logic signed [7:0] weight_0 = 1;
  parameter logic signed [7:0] weight_1 = 2;
  parameter logic signed [7:0] weight_2 = 3;
  parameter logic signed [7:0] weight_3 = 4;

endpackage