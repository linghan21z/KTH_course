package state_pkg;
  typedef enum logic [1:0] {idle = 2'b00, c0 = 2'b01, c1=2'b10 } state_ty;
endpackage