class random_pkg #(parameter N=4);
  rand logic [N-1] a,b;
endclass