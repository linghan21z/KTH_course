library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.types.all;

entity Sigmoid is

	port ( 
		result_in : in signed(INT_BITS+FRAC_BITS-1 downto 0); 
		output    : out signed(INT_BITS+FRAC_BITS-1 downto 0));

end Sigmoid;

architecture Behavioral of Sigmoid is
	-- signal output_tmp : unsigned(INT_BITS+FRAC_BITS-1 downto 0);
Begin
	with result_in select output <= 
		"00000001" when "10000000",
		"00000001" when "10000001",
		"00000001" when "10000010",
		"00000001" when "10000011",
		"00000001" when "10000100",
		"00000001" when "10000101",
		"00000001" when "10000110",
		"00000001" when "10000111",
		"00000001" when "10001000",
		"00000001" when "10001001",
		"00000001" when "10001010",
		"00000001" when "10001011",
		"00000001" when "10001100",
		"00000001" when "10001101",
		"00000001" when "10001110",
		"00000001" when "10001111",
		"00000001" when "10010000",
		"00000001" when "10010001",
		"00000001" when "10010010",
		"00000001" when "10010011",
		"00000001" when "10010100",
		"00000001" when "10010101",
		"00000001" when "10010110",
		"00000001" when "10010111",
		"00000001" when "10011000",
		"00000001" when "10011001",
		"00000001" when "10011010",
		"00000001" when "10011011",
		"00000001" when "10011100",
		"00000001" when "10011101",
		"00000001" when "10011110",
		"00000001" when "10011111",
		"00000010" when "10100000",
		"00000010" when "10100001",
		"00000010" when "10100010",
		"00000010" when "10100011",
		"00000010" when "10100100",
		"00000010" when "10100101",
		"00000010" when "10100110",
		"00000010" when "10100111",
		"00000010" when "10101000",
		"00000010" when "10101001",
		"00000010" when "10101010",
		"00000010" when "10101011",
		"00000010" when "10101100",
		"00000010" when "10101101",
		"00000010" when "10101110",
		"00000010" when "10101111",
		"00000010" when "10110000",
		"00000010" when "10110001",
		"00000011" when "10110010",
		"00000011" when "10110011",
		"00000011" when "10110100",
		"00000011" when "10110101",
		"00000011" when "10110110",
		"00000011" when "10110111",
		"00000011" when "10111000",
		"00000011" when "10111001",
		"00000011" when "10111010",
		"00000011" when "10111011",
		"00000011" when "10111100",
		"00000100" when "10111101",
		"00000100" when "10111110",
		"00000100" when "10111111",
		"00000100" when "11000000",
		"00000100" when "11000001",
		"00000100" when "11000010",
		"00000100" when "11000011",
		"00000100" when "11000100",
		"00000100" when "11000101",
		"00000100" when "11000110",
		"00000101" when "11000111",
		"00000101" when "11001000",
		"00000101" when "11001001",
		"00000101" when "11001010",
		"00000101" when "11001011",
		"00000101" when "11001100",
		"00000101" when "11001101",
		"00000110" when "11001110",
		"00000110" when "11001111",
		"00000110" when "11010000",
		"00000110" when "11010001",
		"00000110" when "11010010",
		"00000110" when "11010011",
		"00000110" when "11010100",
		"00000111" when "11010101",
		"00000111" when "11010110",
		"00000111" when "11010111",
		"00000111" when "11011000",
		"00000111" when "11011001",
		"00000111" when "11011010",
		"00001000" when "11011011",
		"00001000" when "11011100",
		"00001000" when "11011101",
		"00001000" when "11011110",
		"00001000" when "11011111",
		"00001001" when "11100000",
		"00001001" when "11100001",
		"00001001" when "11100010",
		"00001001" when "11100011",
		"00001001" when "11100100",
		"00001010" when "11100101",
		"00001010" when "11100110",
		"00001010" when "11100111",
		"00001010" when "11101000",
		"00001010" when "11101001",
		"00001011" when "11101010",
		"00001011" when "11101011",
		"00001011" when "11101100",
		"00001011" when "11101101",
		"00001100" when "11101110",
		"00001100" when "11101111",
		"00001100" when "11110000",
		"00001100" when "11110001",
		"00001101" when "11110010",
		"00001101" when "11110011",
		"00001101" when "11110100",
		"00001101" when "11110101",
		"00001110" when "11110110",
		"00001110" when "11110111",
		"00001110" when "11111000",
		"00001110" when "11111001",
		"00001111" when "11111010",
		"00001111" when "11111011",
		"00001111" when "11111100",
		"00001111" when "11111101",
		"00010000" when "11111110",
		"00010000" when "11111111",
		"00010000" when "00000000",
		"00010000" when "00000001",
		"00010000" when "00000010",
		"00010001" when "00000011",
		"00010001" when "00000100",
		"00010001" when "00000101",
		"00010001" when "00000110",
		"00010010" when "00000111",
		"00010010" when "00001000",
		"00010010" when "00001001",
		"00010010" when "00001010",
		"00010011" when "00001011",
		"00010011" when "00001100",
		"00010011" when "00001101",
		"00010011" when "00001110",
		"00010100" when "00001111",
		"00010100" when "00010000",
		"00010100" when "00010001",
		"00010100" when "00010010",
		"00010101" when "00010011",
		"00010101" when "00010100",
		"00010101" when "00010101",
		"00010101" when "00010110",
		"00010110" when "00010111",
		"00010110" when "00011000",
		"00010110" when "00011001",
		"00010110" when "00011010",
		"00010110" when "00011011",
		"00010111" when "00011100",
		"00010111" when "00011101",
		"00010111" when "00011110",
		"00010111" when "00011111",
		"00010111" when "00100000",
		"00011000" when "00100001",
		"00011000" when "00100010",
		"00011000" when "00100011",
		"00011000" when "00100100",
		"00011000" when "00100101",
		"00011001" when "00100110",
		"00011001" when "00100111",
		"00011001" when "00101000",
		"00011001" when "00101001",
		"00011001" when "00101010",
		"00011001" when "00101011",
		"00011010" when "00101100",
		"00011010" when "00101101",
		"00011010" when "00101110",
		"00011010" when "00101111",
		"00011010" when "00110000",
		"00011010" when "00110001",
		"00011010" when "00110010",
		"00011011" when "00110011",
		"00011011" when "00110100",
		"00011011" when "00110101",
		"00011011" when "00110110",
		"00011011" when "00110111",
		"00011011" when "00111000",
		"00011011" when "00111001",
		"00011100" when "00111010",
		"00011100" when "00111011",
		"00011100" when "00111100",
		"00011100" when "00111101",
		"00011100" when "00111110",
		"00011100" when "00111111",
		"00011100" when "01000000",
		"00011100" when "01000001",
		"00011100" when "01000010",
		"00011100" when "01000011",
		"00011101" when "01000100",
		"00011101" when "01000101",
		"00011101" when "01000110",
		"00011101" when "01000111",
		"00011101" when "01001000",
		"00011101" when "01001001",
		"00011101" when "01001010",
		"00011101" when "01001011",
		"00011101" when "01001100",
		"00011101" when "01001101",
		"00011101" when "01001110",
		"00011110" when "01001111",
		"00011110" when "01010000",
		"00011110" when "01010001",
		"00011110" when "01010010",
		"00011110" when "01010011",
		"00011110" when "01010100",
		"00011110" when "01010101",
		"00011110" when "01010110",
		"00011110" when "01010111",
		"00011110" when "01011000",
		"00011110" when "01011001",
		"00011110" when "01011010",
		"00011110" when "01011011",
		"00011110" when "01011100",
		"00011110" when "01011101",
		"00011110" when "01011110",
		"00011110" when "01011111",
		"00011110" when "01100000",
		"00011111" when "01100001",
		"00011111" when "01100010",
		"00011111" when "01100011",
		"00011111" when "01100100",
		"00011111" when "01100101",
		"00011111" when "01100110",
		"00011111" when "01100111",
		"00011111" when "01101000",
		"00011111" when "01101001",
		"00011111" when "01101010",
		"00011111" when "01101011",
		"00011111" when "01101100",
		"00011111" when "01101101",
		"00011111" when "01101110",
		"00011111" when "01101111",
		"00011111" when "01110000",
		"00011111" when "01110001",
		"00011111" when "01110010",
		"00011111" when "01110011",
		"00011111" when "01110100",
		"00011111" when "01110101",
		"00011111" when "01110110",
		"00011111" when "01110111",
		"00011111" when "01111000",
		"00011111" when "01111001",
		"00011111" when "01111010",
		"00011111" when "01111011",
		"00011111" when "01111100",
		"00011111" when "01111101",
		"00011111" when "01111110",
		"00011111" when "01111111",
		"00000000" when others; 
	-- output <= to_sfixed(unsigned(output_tmp), INT_BITS, -FRAC_BITS);
end Behavioral;
	
